`timescale 1 ns/100 ps

module reg_4bit ( input ld,
                  input clk,
                  input [0:3] d,
                  output [0:3] q);
// Inserir codigo para funcionamento do registrador de 4 bits.
endmodule
