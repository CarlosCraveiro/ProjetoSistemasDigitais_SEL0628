`timescale 1 ns/100 ps

module counter_block( input enable,
                      input reset,
                      input clk,
                      input load,
                      output [0:6] ssg,
                      output enable_next);
// Implementar logica de funcionamento do bloco de contagem
endmodule
