`timescale 1 ns/100 ps

module d_slp_counter( input enable,
                      input reset,
                      input load,
                      output [6:0] ssg_1,
                      output [6:0] ssg_2,
                      output [6:0] ssg_3, 
                      output en_machine);
// Implementar funcionamento do contador presente no ADC de Rampa Dupla
endmodule

