`timescale 1 ns/100 ps

module counter_bcd(  input clk,
                        input enable,
                        input reset,
                        output reg [0:3] bcd,
                        output cnt_9);
// Implementar funcionamento do modulo contador BCD
endmodule
