`timescale 1 ns/100 ps

module bcd_to_ssg ( input [3:0] bcd,
                    output [6:0] ssg);
// Inserir codigo de funcionamento para conversor bcd para sete segmentos
endmodule
