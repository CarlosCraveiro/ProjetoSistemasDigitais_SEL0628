`timescale 1 ns/100 ps

module control_machine( input start,
                        input clk,
                        input finished_counting,
                        input cap_discharged,
                        output ch_Vmeasured,
                        output ch_Vref,
                        output ch_Zero,
                        output reset,
                        output enable_counting);
  // Implementar logica de controle de ADC do tipo rampa dupla
endmodule
