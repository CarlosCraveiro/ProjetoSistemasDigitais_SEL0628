`timescale 1 ns/100 ps

module bcd_to_ssg ( input [0:3] bcd,
                    output [0:6] ssg);
// Inserir codigo de funcionamento para conversor bcd para sete segmentos
endmodule
