`timescale 1 ns/100 ps

module d_slp_counter( input enable,
                      input reset,
                      input load,
                      output [0:6] ssg_1,
                      output [0:6] ssg_2,
                      output [0:6] ssg_3, 
                      output en_machine);
// Implementar funcionamento do contador presente no ADC de Rampa Dupla
endmodule

